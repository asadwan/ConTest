contextModel TranslationApp {	
	
	// Mark: context declaration 
	
	context INTERNET_CONNECTIVITY {
		providers: [WIFI_ADAPTER, CELL_ADAPTER],
		properties: [connectivity: Connectivity],
	}
	
	context LOCATION {
		providers: [GPS_SENSOR, CELL_ADAPTER],
		properties: [availability: Availability, longitude: double, latitude: double],
	}
	
	context COUNTRY derives LOCATION {
		properties: [country: Country],
		mappings: {
			country.france -> LOCATION.longitude == "x" and LOCATION.latitude == "y", // a specific value or range of values 
			country.germany -> LOCATION.longitude == "x" and LOCATION.latitude == "y",
			country.spain -> LOCATION.longitude == "x" and LOCATION.latitude == "y"
		}
	}
	
	static context OS {
		providers: [DEVICE_API],
		properties: [os: OS],
	}
	
	static context SCREEN_ORIENTATION {
		providers: [GYROSCOPE_SENSOR],
		properties: [orientation: Screen_Orientation],
	}
	
	// Mark: context providers declaration
	
	providers {
		WIFI_ADAPTER,
		CELL_ADAPTER,
		GPS_SENSOR,
		DEVICE_API,
		GYROSCOPE_SENSOR
	}	
	
	// Mark: situations declaration
	
	
	situation INTERNET_DISCONNECTED {
		INTERNET_CONNECTIVITY.connectivity == offline
	}
	
	
	situation LOCATION_UNAVAILABLE {
		LOCATION.availability == unavailable
	}
	
	// Mark: context data types declaration
	
	type Connectivity {offline, wifi, slow3G, fast3G, _4g, high_latency}
	
	type OS {android, ios}
	
	type Screen_Orientation {portrait, landscape}
	
	type Country {france, germany, spain, uk}
	
	type Availability {available, unavailable}
	
}